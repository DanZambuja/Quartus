library IEEE;
use IEEE.std_logic_1164.all;

entity deMux_4 is
	port (SEL : in std_logic_vector(3 downto 0);
			E: in std_logic_vector(15 downto 0);
			S1, S2, S3, S4: out std_logic_vector(15 downto 0));

end deMux_4;


architecture behavioral of deMux_4 is
begin
process(SEL)
begin
	if (SEL = "0001") then
		S1 <= E;
	elsif (SEL = "0010") then
		S2 <= E;
	elsif (SEL = "0011") then 
		S3 <= E;
	elsif (SEL = "0100") then 
		S4 <= E;
	end if;
end process;
end behavioral;