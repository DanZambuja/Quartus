library IEEE;
use IEEE.std_logic_1164.all;

entity contador2bits is 

	port (clock, reset, enable: in std_logic;
			saida: out std_logic_vector(1 downto 0));
	
end contador2bits;


architecture arch of contador2bits is


begin




end arch;